module sim_top
    (
        input clk,
        input rst,
        inout sio3
    );

endmodule

