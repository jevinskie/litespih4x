module TristateModelHand
    (
        input clk,
        input rst,
        inout SIO3
    );

    assign SIO3 = 1'b0;

endmodule

