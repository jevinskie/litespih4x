module sim_top
    (
        input sys_clk,
        input sys_rst,
        inout sio3
    );

endmodule

