module TristateModelHand
    (
        input clk,
        input rst,
        inout sio3
    );

    assign sio3 = 1'b0;

endmodule

